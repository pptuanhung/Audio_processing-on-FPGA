package Genwave_Pkg; // PACKAGE

  parameter int GEN_WD = 16;
  parameter int DC_WD  = 4;
  parameter int N_WD   = 16;

endpackage: Genwave_Pkg
