module data_out 
