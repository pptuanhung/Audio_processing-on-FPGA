module show_led_4 (
  input  logic  [1:0] sel,
  output logic  [6:0] out
);
  always@(*)  begin
    case(sel)
        2'b00: out <= 7'b0010010; //S 
        2'b01: out <= 7'b1001000; //n
        2'b10: out <= 7'b1000010; //G
        2'b11: out <= 7'b1111111; //no

    endcase
  end
endmodule