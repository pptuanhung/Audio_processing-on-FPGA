module core 


//data_in



// control 



//data_process



//data_out


endmodule